
module add_32()






endmodule