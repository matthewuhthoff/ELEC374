
module alu(
    input clk, clear, incrementPC, branch

    input wire[31:0] a_reg,
    
)




endmodule